`ifndef MACROS_SV
`define MACROS_SV

`define REGBITS  5
`define OPFUNC  10
`define IMMREG  12
`define INSTRSZ 32

`endif
