typedef enum {
    reg_zero = 5'b00000,
    reg_ra = 5'b00001,
    reg_sp = 5'b00010,
    reg_gp = 5'b00011,
    reg_tp = 5'b00100,
    reg_t0 = 5'b00101,
    reg_t1 = 5'b00110,
    reg_t2 = 5'b00111,
    reg_s0 = 5'b01000,
    reg_s1 = 5'b01001,
    reg_a0 = 5'b01010,
    reg_a1 = 5'b01011,
    reg_a2 = 5'b01100,
    reg_a3 = 5'b01101,
    reg_a4 = 5'b01110,
    reg_a5 = 5'b01111,
    reg_a6 = 5'b10000,
    reg_a7 = 5'b10001,
    reg_s2 = 5'b10010,
    reg_s3 = 5'b10011,
    reg_s4 = 5'b10100,
    reg_s5 = 5'b10101,
    reg_s6 = 5'b10110,
    reg_s7 = 5'b10111,
    reg_s8 = 5'b11000,
    reg_s9 = 5'b11001,
    reg_s10 = 5'b11010,
    reg_s11 = 5'b11011,
    reg_t3 = 5'b11100,
    reg_t4 = 5'b11101,
    reg_t5 = 5'b11110,
    reg_t6 = 5'b11111
} register_enum;

logic [63:0] register_file[31:0];
