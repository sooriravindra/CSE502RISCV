typedef enum {INITIAL, WAIT_RESP, GOT_RESP} State;
State state, next_state;
